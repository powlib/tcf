`timescale 1ns / 1ps

module test_ipmaxi();

  initial begin
    $dumpfile("waveform.vcd");
    //$dumpvars(10, dut0);
  end  

endmodule